// Optimized via extended random search (150 trials)
// Accuracy: 75.0%

parameter WEIGHT_I0_H0 = 15;
parameter WEIGHT_I0_H1 = 0;
parameter WEIGHT_I0_H2 = 0;
parameter WEIGHT_I0_H3 = 0;
parameter WEIGHT_I0_H4 = 8;
parameter WEIGHT_I0_H5 = 0;
parameter WEIGHT_I0_H6 = 8;
parameter WEIGHT_I0_H7 = 0;
parameter WEIGHT_I1_H0 = 0;
parameter WEIGHT_I1_H1 = 15;
parameter WEIGHT_I1_H2 = 0;
parameter WEIGHT_I1_H3 = 0;
parameter WEIGHT_I1_H4 = 8;
parameter WEIGHT_I1_H5 = 0;
parameter WEIGHT_I1_H6 = 0;
parameter WEIGHT_I1_H7 = 8;
parameter WEIGHT_I2_H0 = 0;
parameter WEIGHT_I2_H1 = 0;
parameter WEIGHT_I2_H2 = 15;
parameter WEIGHT_I2_H3 = 0;
parameter WEIGHT_I2_H4 = 0;
parameter WEIGHT_I2_H5 = 8;
parameter WEIGHT_I2_H6 = 8;
parameter WEIGHT_I2_H7 = 0;
parameter WEIGHT_I3_H0 = 0;
parameter WEIGHT_I3_H1 = 0;
parameter WEIGHT_I3_H2 = 0;
parameter WEIGHT_I3_H3 = 15;
parameter WEIGHT_I3_H4 = 0;
parameter WEIGHT_I3_H5 = 8;
parameter WEIGHT_I3_H6 = 0;
parameter WEIGHT_I3_H7 = 8;

parameter WEIGHT_H0_O0 = 0;
parameter WEIGHT_H0_O1 = 0;
parameter WEIGHT_H0_O2 = 0;
parameter WEIGHT_H1_O0 = 0;
parameter WEIGHT_H1_O1 = 0;
parameter WEIGHT_H1_O2 = 0;
parameter WEIGHT_H2_O0 = 1;
parameter WEIGHT_H2_O1 = 0;
parameter WEIGHT_H2_O2 = 3;
parameter WEIGHT_H3_O0 = 0;
parameter WEIGHT_H3_O1 = 0;
parameter WEIGHT_H3_O2 = 2;
parameter WEIGHT_H4_O0 = 0;
parameter WEIGHT_H4_O1 = 15;
parameter WEIGHT_H4_O2 = 0;
parameter WEIGHT_H5_O0 = 15;
parameter WEIGHT_H5_O1 = 3;
parameter WEIGHT_H5_O2 = 15;
parameter WEIGHT_H6_O0 = 15;
parameter WEIGHT_H6_O1 = 0;
parameter WEIGHT_H6_O2 = 0;
parameter WEIGHT_H7_O0 = 0;
parameter WEIGHT_H7_O1 = 15;
parameter WEIGHT_H7_O2 = 15;

parameter BIAS_OUTPUT_0 = 0;
parameter BIAS_OUTPUT_1 = 0;
parameter BIAS_OUTPUT_2 = 0;
